module MuxH (
input wire[31:0] FromB,
input wire[31:0] Immediate,
input wire[0:0] ShiftAmt,
output reg[31:0] toShift
);
parameter S0 = 0, S1 = 1;
always @(*) begin
	case(ShiftAmt)
		S0:
			toShift <= FromB;
		S1:
			toShift <= Immediate;
	endcase
end

endmodule