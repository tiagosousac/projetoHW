module CPU (clock, reset, AluResult, MuxIOut, MuxFOut, MuxGOut, MuxHOut, AluOp, RegAOut, RegBOut, RegPCOut, MemData, estado);

input clock;
input reset;

output reg [31:0] AluResult;
wire [31:0] SSOut, RegWriteOutA, RegWriteOutB, MuxEOut, RegEPCOut, RegAluOutOut,  RegMDROut;
wire [31:0] HICtrlOut, RegHIOut, LOCtrlOut, RegLOOut, RegDeslocOut, MuxCOut, MuxDOut, Extend16a32Out, OffsetExtendidoLeft2;
wire [4:0] RS, RT, RD, MuxBOut;
wire [15:0] Offset;
wire [5:0] Opcode;
output wire [31:0] RegAOut, RegBOut, RegPCOut, MemData;
output wire [6:0] estado;
wire [5:0] Funct;
output wire [31:0] MuxIOut;
output wire [31:0] MuxFOut;
output wire [31:0] MuxGOut;
output wire [31:0] MuxHOut;

wire [4:0] BCut, Shamt;
assign BCut = RegBOut[4:0];
assign Shamt = Offset[10:6];
assign RD = Offset[15:11];

wire MuxAOut;
wire WriteCond;
wire PCWrite;
wire RegWrite;
wire Wr;
wire IRWrite;
wire WriteRegA;
wire WriteRegB;
wire AluOutControl;
wire EPCWrite;
wire ShiftSrc;
wire ShiftAmt;
wire DivCtrl;
wire MultCtrl;
wire HICtrl;
wire LOCtrl;
wire WriteHI;
wire WriteLO;
wire MDRCtrl;
wire [1:0] ExceptionCtrl;

wire [1:0] AluSrcA;
wire [2:0] AluSrcB;
output wire [2:0] AluOp;
wire [2:0] PCSource;
wire [2:0] IorD;
wire [2:0] ShiftCtrl;
wire [2:0] RegDst;
wire [3:0] MemToReg;

Registrador registradorA(clock, reset, WriteRegA, RegWriteOutA, RegAOut);
Registrador registradorB(clock, reset, WriteRegB, RegWriteOutB, RegBOut);
Registrador PC (clock, reset, PCWrite, MuxEOut, RegPCOut);
Registrador EPC (clock, reset, EPCWrite, AluOut, RegEPCOut);
Registrador AluOut (clock, reset, AluOutControl, AluResult, RegAluOutOut);
Registrador MDR(clock, reset, MDRCtrl, MemData, RegMDROut);
Registrador HI(clock, reset, WriteHI, HICtrlOut, RegHIOut);
Registrador LO(clock, reset, WriteLO, LOCtrlOut, RegLOOut);
Banco_reg banco_registradores(clock, reset, RegWrite, RS, RT, MuxBOut, MuxIOut, RegWriteOutA, RegWriteOutB);
RegDesloc regdesloc(clock, reset, ShiftCtrl, MuxHOut, MuxGOut, RegDeslocOut);
Controle controle(clock, reset, Opcode, Funct, WriteCond,PCWrite,RegWrite,Wr,IRWrite,WriteRegA,WriteRegB,AluOutControl,EPCWrite,ShiftSrc,ShiftAmt,DivCtrl,MultCtrl,HICtrl,LOCtrl,WriteHI,WriteLO,MDRCtrl,ExceptionCtrl, AluSrcA,AluSrcB,AluOp,PCSource,IorD,ShiftCtrl,RegDst,MemToReg, estado);
Memoria memoria(MuxAOut, clock, Wr, SSOut, MemData);
Instr_Reg InstructionRegisters (clock, reset, IRWrite, MemData, Opcode, RS, RT, Offset);	
ula32 Alu(MuxCOut, MuxDOut, AluOp, AluResult, Overflow, Negativo, Zero, EQ, GT, LT);

//Declara�ao de cada Mux
MuxA MuxA(RegPCOut, MuxFOut, AluResult, RegAluOutOut, RegAOut, IorD, MuxAOut);
MuxB MuxB(RS, RT, RD, RegDst, MuxBOut);
MuxC MuxC(RegPCOut, RegBOut, RegAOut, MemData, AluSrcA, MuxCOut);
MuxD MuxD(RegBOut, Extend16a32Out, RegMDROut, OffsetExtendidoLeft2, AluSrcB, MuxDOut);
MuxE MuxE(RegAOut, AluResult, 1'd0, RegAluOutOut, RegEPCOut, 1'd0, PCSource, MuxEOut);
MuxF MuxF(ExceptionCtrl, MuxFOut);
MuxG MuxG(RegAOut, RegBOut, ShiftSrc, MuxGOut);
MuxH MuxH(BCut, Shamt, ShiftAmt, MuxHOut); //Mudar nome Bcut
MuxI MuxI(LT, LoadOut, RegDeslocOut, RegHIOut, RegLOOut, RegBOut, RegAOut, RegAluOutOut, OffsetExtendidoLeft2, OffsetExtendidoLeft16, MemToReg, MuxIOut); //LoadOut = saida da caixa Load apos MDR; OffsetExtendidoLeft16 = saida do shift left 16, acredito que ainda nao inicializada

SE1632 SignExtend16a32(Offset, OffsetExtendido);
ShiftLeft2 sl2(OffsetExtendido, OffsetExtendidoLeft2);
FunctExtract functextract(Offset, Funct);


endmodule